LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY Group_3 IS
PORT ( CLK50MHZ : IN  STD_LOGIC;
		 KEY      : IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		 SW       : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		 LEDR     : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		 HEX0     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX1     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX2     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX3     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX4     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 HEX5     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 GPIO     : OUT STD_LOGIC_VECTOR(36 DOWNTO 0)
		 );
END ENTITY Group_3;


ARCHITECTURE behaviour OF Group_3 IS
SIGNAL CLK_play         : STD_LOGIC;
SIGNAL CLK_ALM          : STD_LOGIC;
SIGNAL BUZZ             : STD_LOGIC;
SIGNAL RSEST, STRT, STP : STD_LOGIC;
SIGNAL SEC_FLIP_0       : STD_LOGIC:='1';
SIGNAL MIN_FLIP_0       : STD_LOGIC:='1';
SIGNAL K                : STD_LOGIC:='0';
SIGNAL SET              : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL ALARM            : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL ALM_LIGHT        : STD_LOGIC_VECTOR(8 DOWNTO 0);

BEGIN

STRT             <=          KEY(0);
STP              <=          KEY(1);
RSEST            <=           SW(9);
SET              <=  SW(1 DOWNTO 0);

GPIO(5)          <=            BUZZ;
LEDR(9)          <=               K;
LEDR(8 DOWNTO 0) <=       ALM_LIGHT;

DISP_CLK_3: WORK.Pl_CLK  PORT MAP(clk_3 => CLK50MHZ,
											T2     => CLK_play);
DISP_CLK_4: WORK.ALM_CLK PORT MAP(clk_4 => CLK50MHZ,
											T3     => CLK_ALM);

PROCESS(CLK_play, RSEST, SEC_FLIP_0, MIN_FLIP_0, STRT, STP, K, BUZZ)

VARIABLE P1_0, P2_0, P3_0 : INTEGER := 0;
VARIABLE P2_1_0, P3_1_0   : INTEGER := 0;
VARIABLE ALM_H, ALM_M     : INTEGER := 0;
BEGIN

IF SET = "00" THEN
		
		IF RISING_EDGE(STRT) THEN
			IF RSEST = '0' THEN
				ALM_M := 0;
			ELSE
				IF ALM_M = 59 THEN
					ALM_M := 0;
				ELSE
					ALM_M := ALM_M + 1;
				END IF;
			END IF;
		END IF;
		
		IF RISING_EDGE(STP) THEN
			IF RSEST = '0' THEN
				ALM_H := 0;
			ELSE
				IF ALM_H = 23 THEN
					ALM_H := 0;
				ELSE
					ALM_H := ALM_H + 1;
				END IF;
			END IF;
		END IF;
		
		P2_0 := ALM_M;
		
		P3_0 := ALM_H;
		
		IF    P2_0 = 0 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 1 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 2 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 3 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 4 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 5 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 6 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 7 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 8 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 9 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 10 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 11 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 12 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 13 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 14 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 15 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 16 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 17 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 18 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 19 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 20 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 21 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 22 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 23 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 24 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 25 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 26 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 27 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 28 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 29 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 30 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 31 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 32 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 33 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 34 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 35 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 36 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 37 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 38 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 39 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 40 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 41 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 42 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 43 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 44 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 45 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 46 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 47 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 48 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 49 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 50 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 51 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 52 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 53 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 54 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 55 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 56 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 57 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 58 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 59 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSE
			HEX2 <= STD_LOGIC_VECTOR'("01111111");
			HEX3 <= STD_LOGIC_VECTOR'("01111111");
		END IF;
		
		IF P3_0 = 0 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 1 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 2 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 3 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 4 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 5 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 6 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 7 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 8 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 9 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 10 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 11 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 12 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 13 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 14 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 15 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 16 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 17 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 18 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 19 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 20 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 21 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 22 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 23 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSE
			HEX4 <= STD_LOGIC_VECTOR'("01111111");
			HEX5 <= STD_LOGIC_VECTOR'("01111111");
		END IF;
		
	
	ELSIF SET = "01" THEN
		
		IF RISING_EDGE(STRT) THEN
			IF RSEST = '0' THEN
				P2_1_0 := 0;
			ELSE
				IF P2_1_0 = 59 THEN
					P2_1_0 := 0;
				ELSE
					P2_1_0 := P2_1_0 + 1;
				END IF;
			END IF;
		END IF;
		
		IF RISING_EDGE(STP) THEN
			IF RSEST = '0' THEN
				P3_1_0 := 0;
			ELSE
				IF P3_1_0 = 23 THEN
					P3_1_0 := 0;
				ELSE
					P3_1_0 := P3_1_0 + 1;
				END IF;
			END IF;
		END IF;
		
		P2_0 := P2_1_0;
		
		P3_0 := P3_1_0;
		
		IF    P2_0 = 0 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 1 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 2 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 3 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 4 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 5 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 6 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 7 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 8 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 9 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 10 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 11 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 12 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 13 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 14 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 15 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 16 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 17 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 18 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 19 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 20 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 21 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 22 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 23 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 24 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 25 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 26 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 27 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 28 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 29 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 30 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 31 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 32 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 33 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 34 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 35 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 36 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 37 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 38 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 39 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 40 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 41 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 42 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 43 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 44 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 45 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 46 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 47 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 48 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 49 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 50 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 51 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 52 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 53 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 54 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 55 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 56 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 57 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 58 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 59 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSE
			HEX2 <= STD_LOGIC_VECTOR'("01111111");
			HEX3 <= STD_LOGIC_VECTOR'("01111111");
		END IF;
		
		IF P3_0 = 0 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 1 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 2 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 3 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 4 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 5 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 6 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 7 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 8 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 9 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 10 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 11 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 12 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 13 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 14 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 15 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 16 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 17 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 18 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 19 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 20 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 21 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 22 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 23 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSE
			HEX4 <= STD_LOGIC_VECTOR'("01111111");
			HEX5 <= STD_LOGIC_VECTOR'("01111111");
		END IF;
		
	ELSE
		
		IF (P3_0 = ALM_H) AND (P2_0 = ALM_M) THEN
			IF SW(8) = '0' THEN
				K <= '1';
				BUZZ <= '1';
				IF RISING_EDGE(CLK_ALM) THEN
					ALM_LIGHT <= NOT(ALM_LIGHT);
				END IF;
			ELSE
				K <= '0';
				BUZZ <= '0';
			END IF;
		ELSE
			K <= '0';
			BUZZ <= '0';
		END IF;
		
		IF RISING_EDGE(CLK_play) THEN
					
			IF RSEST = '1' THEN
				P1_0 := P1_0 + 1;
			ELSE
				P1_0 := 0;
			END IF;
			
			IF (P1_0 = 60) THEN
				SEC_FLIP_0 <= '0';
				P1_0 :=   0;
			ELSE
				SEC_FLIP_0 <= '1';
				P1_0 :=   P1_0;
			END IF;
			
			IF P1_0 = 0 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 1 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 2 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 3 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 4 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 5 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 6 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 7 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 8 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 9 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("11000000");
			ELSIF P1_0 = 10 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 11 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 12 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 13 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 14 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 15 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 16 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 17 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 18 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 19 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("11111001");
			ELSIF P1_0 = 20 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 21 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 22 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 23 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 24 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 25 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 26 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 27 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 28 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 29 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10100100");
			ELSIF P1_0 = 30 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 31 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 32 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 33 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 34 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 35 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 36 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 37 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 38 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 39 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10110000");
			ELSIF P1_0 = 40 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 41 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 42 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 43 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 44 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 45 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 46 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 47 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 48 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 49 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10011001");
			ELSIF P1_0 = 50 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01000000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 51 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111001");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 52 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00100100");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 53 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00110000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 54 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011001");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 55 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00010010");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 56 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000010");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 57 THEN
				HEX0 <= STD_LOGIC_VECTOR'("01111000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 58 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00000000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSIF P1_0 = 59 THEN
				HEX0 <= STD_LOGIC_VECTOR'("00011000");
				HEX1 <= STD_LOGIC_VECTOR'("10010010");
			ELSE
				HEX0 <= STD_LOGIC_VECTOR'("01111111");
				HEX1 <= STD_LOGIC_VECTOR'("01111111");
			END IF;
				
		END IF;
			
		IF RSEST = '1' THEN
			IF FALLING_EDGE(SEC_FLIP_0) THEN
				P2_0 := P2_0 + 1;
			END IF;
		ELSE
			P2_0 := 0;
		END IF;
			
		IF (P2_0 = 60) THEN
			MIN_FLIP_0 <= '0';
			P2_0 :=   0;
		ELSE
			MIN_FLIP_0 <= '1';
			P2_0 :=   P2_0;
		END IF;
		
		IF    P2_0 = 0 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 1 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 2 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 3 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 4 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 5 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 6 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 7 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 8 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 9 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P2_0 = 10 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 11 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 12 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 13 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 14 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 15 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 16 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 17 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 18 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 19 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P2_0 = 20 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 21 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 22 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 23 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 24 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 25 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 26 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 27 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 28 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 29 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P2_0 = 30 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 31 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 32 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 33 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 34 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 35 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 36 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 37 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 38 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 39 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10110000");
		ELSIF P2_0 = 40 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 41 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 42 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 43 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 44 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 45 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 46 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 47 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 48 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 49 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10011001");
		ELSIF P2_0 = 50 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 51 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 52 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00100100");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 53 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00110000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 54 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011001");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 55 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00010010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 56 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000010");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 57 THEN
			HEX2 <= STD_LOGIC_VECTOR'("01111000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 58 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00000000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSIF P2_0 = 59 THEN
			HEX2 <= STD_LOGIC_VECTOR'("00011000");
			HEX3 <= STD_LOGIC_VECTOR'("10010010");
		ELSE
			HEX2 <= STD_LOGIC_VECTOR'("01111111");
			HEX3 <= STD_LOGIC_VECTOR'("01111111");
		END IF;
		
		IF RSEST = '1' THEN
			IF FALLING_EDGE(MIN_FLIP_0) THEN
				P3_0 := P3_0 + 1;
			END IF;
		ELSE
			P3_0 := 0;
		END IF;
		
		IF (P3_0 = 24) THEN
			P3_0 := 0;
		ELSE
			P3_0 := P3_0;
		END IF;
		
		IF P3_0 = 0 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 1 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 2 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 3 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 4 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 5 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 6 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 7 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 8 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 9 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11000000");
		ELSIF P3_0 = 10 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 11 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 12 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 13 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 14 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011001");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 15 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00010010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 16 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000010");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 17 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 18 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00000000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 19 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00011000");
			HEX5 <= STD_LOGIC_VECTOR'("11111001");
		ELSIF P3_0 = 20 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01000000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 21 THEN
			HEX4 <= STD_LOGIC_VECTOR'("01111001");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 22 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00100100");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSIF P3_0 = 23 THEN
			HEX4 <= STD_LOGIC_VECTOR'("00110000");
			HEX5 <= STD_LOGIC_VECTOR'("10100100");
		ELSE
			HEX4 <= STD_LOGIC_VECTOR'("01111111");
			HEX5 <= STD_LOGIC_VECTOR'("01111111");
		END IF;
			
	END IF;
	
END PROCESS;
END behaviour;